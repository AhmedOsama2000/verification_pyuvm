package alu_pkg;
	
	`include "transaction.sv"
	`include "driver.sv"
	`include "monitor.sv"
	`include "sequencer.sv"
	`include "env.sv"

endpackage